package uvm_tb_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "../uvm_tb/my_item.sv"
    `include "../uvm_tb/my_sequence.sv"
    `include "../uvm_tb/my_sequencer.sv"
    `include "../uvm_tb/my_driver.sv"
    `include "../uvm_tb/my_monitor.sv"
    `include "../uvm_tb/my_agent.sv"
    `include "../uvm_tb/my_scoreboard.sv"
    `include "../uvm_tb/my_env.sv"
    `include "../uvm_tb/my_test.sv"



endpackage : uvm_tb_pkg
