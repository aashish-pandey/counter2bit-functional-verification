interface counter_if;
    logic clk;
    logic reset;
    logic up_down;
    logic [1:0] count;
endinterface